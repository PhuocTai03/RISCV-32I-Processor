`timescale 1ns / 1ps
module StallingUnit(

    );
    
    
endmodule